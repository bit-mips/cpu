`ifndef MIPS32R2_CP0_SVH
`define MIPS32R2_CP0_SVH

`define CP0_OPT_ARCH_REV_REL1 0
`define CP0_OPT_ARCH_REV_REL2 1

`define CP0_CMD_READREG  0
/* Read CP0 registers
* no: Reg No
* sel: Reg Sel
* resp: Reg content
*/
`define CP0_CMD_WRITEREG 1
/* Write to CP0 registers
* no: Reg No
* sel: Reg Sel
* data: Write data
*/
`define CP0_CMD_DI       2
/* Disable interrupt
* resp: Status content
*/
`define CP0_CMD_EI       3
/* Enable interrupt */
`define CP0_CMD_TLBPROBE 4
/* TLB Probe */
`define CP0_CMD_TLBREAD  5
/* TLB Read */
`define CP0_CMD_TLBWI    6
/* TLB Write Indexed
* resp: 0 - ok, 1 - CpU, 2 - MCheck
*/
`define CP0_CMD_TLBWR    7
/* TLB Write Random
* resp: 0 - ok, 1 - CpU, 2 - MCheck
*/
`define CP0_CMD_CINVL    8
/* Invalidate all cache data */
`define CP0_CMD_CSYNC    9
/* Writeback all dirty data */
`define CP0_CMD_CHKPRIV  10
/* Check kernel privilege
* resp: 0 - currently in kernel mode, 1 - in user mode
*/

/* Exception generated by CP0 */
/* HardReset */
/* SoftReset */
/* NMI */
`define CP0_EX_INTERRUPT /* external interrupts */          6'h00 /* Int */
`define CP0_EX_MACHCHK /* machine check */                  6'h18 /* MCheck */

/* Exception generated by execution units */
`define CP0_EX_MEM_WRITE /* writing to a non-dirty page */  6'h01 /* Mod */
/* args:
* a0: failing address
*/
`define CP0_EX_IF_TLBMISS /* TLB miss fetching inst */      6'h02 /* TLBML */
/* args:
* a0: failing address
*/
`define CP0_EX_IF_TLBINV /* TLB invalid on fetch */         6'h22 /* TLBIL */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_TLBML /* TLB miss on load */             6'h02 /* TLBML */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_TLBIL /* TLB invalid on load */          6'h22 /* TLBIL */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_TLBMS /* TLB miss on store */            6'h03 /* TLBMS */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_TLBIS /* TLB invalid on store */         6'h23 /* TLBIS */
/* args:
* a0: failing address
*/
`define CP0_EX_IF_ADDRERR /* address error fetching inst */ 6'h04 /* AdEL */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_AEL /* address error on load */          6'h04 /* AdEL */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_AES /* address error on store */         6'h05 /* AdES */
/* args:
* a0: failing address
*/
`define CP0_EX_IF_BUSERR /* bus error fetching inst */      6'h06 /* IBE */
`define CP0_EX_BUSERR /* bus error */                       6'h07 /* DBE */
`define CP0_EX_SYSCALL /* syscall */                        6'h08 /* Sys */
`define CP0_EX_BREAK /* break */                            6'h09 /* Bp */
`define CP0_EX_RESERVED /* reserved instruction */          6'h0a /* RI */
`define CP0_EX_CPUNUSABLE /* coprocessor unusable */        6'h0b /* CpU */
/* args:
* a0: coprocessor index
*/
`define CP0_EX_OVERFLOW /* arithmetic overflow */           6'h0c /* Ov */
`define CP0_EX_TRAP /* trap */                              6'h0d /* Tr */
`define CP0_EX_FP /* floating-point exception */            6'h0f /* FPE */
`define CP0_EX_IF_TLBRI /* page marked as unreadable */     6'h13 /* TLBRI */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_RI /* page marked as unreadable */       6'h13 /* TLBRI */
/* args:
* a0: failing address
*/
`define CP0_EX_IF_TLBXI /* page marked as not executable */ 6'h14 /* TLBXI */
/* args:
* a0: failing address
*/
`define CP0_EX_MEM_WATCH /* data watchpoint hit */          6'h17 /* WATCH */

/* Special operation treated in the same way as exception */
`define CP0_EX_ERET /* exception return */                  6'h30

`endif
